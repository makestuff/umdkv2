--
-- Copyright (C) 2010 Chris McClelland
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--  
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
library ieee;

use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity MemoryController is
	port(
		clk           : in    std_logic;  -- 100MHz
		reset         : in    std_logic;
		nWait         : in    std_logic;
		memRequest    : in    std_logic;
		readNotWrite  : in    std_logic;
		dataBus       : inout std_logic_vector(15 downto 0);
		addressBus    : out   std_logic_vector(22 downto 0);
		nADV          : out   std_logic;
		nCE           : out   std_logic;
		CRE           : out   std_logic;
		nWE           : out   std_logic;
		nOE           : out   std_logic;
		ramClk        : out   std_logic;
		busy          : out   std_logic;
		mcrAddrInput  : in    std_logic_vector(22 downto 0);
		mcrDataInput  : in    std_logic_vector(15 downto 0);
		mcrDataOutput : out   std_logic_vector(15 downto 0)
	);
end MemoryController;

architecture Behavioural of MemoryController is

	type State is (
		STATE_RESET,
		
		STATE_REQUEST_BCR_WRITE0,  -- Assert nADV, nCE, inWE & CRE, drive BCR_INIT on addressBus
		STATE_REQUEST_BCR_WRITE1,  -- Just in case RAM is already in sync mode, wait for ramClk rising
		STATE_REQUEST_BCR_WRITE2,  -- Deassert nADV to clock in BCR_INIT, keep asserting nCE, inWE & CRE
		STATE_WAIT_BCR_WRITE,      -- 2x INIT states plus 7x this state gives 90ns, which meets tCW>85ns
		STATE_FINISH_BCR_WRITE,    -- READ operation must start on a rising ramClk edge, so insert wait
		                           -- state if necessary
		STATE_PREPARE_READ,
		STATE_REQUEST_READ,
		STATE_WAIT_READ,
		STATE_FINISH_READ,
		
		STATE_PREPARE_WRITE,
		STATE_REQUEST_WRITE,
		STATE_WAIT_WRITE,
		STATE_FINISH_WRITE,
		
		STATE_IDLE
	);
	signal iThisState, iNextState : State;
	signal iThisCount, iNextCount : unsigned(3 downto 0);
	signal iDataInput, iDataOutput : std_logic_vector(15 downto 0);
	signal iThisMCRDataOutput, iNextMCRDataOutput : std_logic_vector(15 downto 0);
	signal inWE : std_logic;
	signal iThisRamClk, iNextRamClk : std_logic;
	constant ADDR_HIZ : std_logic_vector(22 downto 0) := (others=>'1');
	constant DATA_HIZ : std_logic_vector(15 downto 0) := (others=>'1');
	constant INIT_BCR : std_logic_vector(22 downto 0) :=
		  "000"  -- Reserved
		& "10"   -- Select BCR
		& "00"   -- Reserved
		& "0"    -- Synchronous mode
		& "1"    -- Fixed initial latency
		& "011"  -- With four cycles latency, max clock for -70x RAM is 52MHz
		& "0"    -- nWait is active low
		& "0"    -- Reserved
		& "0"    -- Assert nWait during delay (data ready first clock after deasserts)
		& "0"    -- Reserved
		& "0"    -- Reserved
		& "01"   -- 1/2-power drive
		& "1"    -- Burst no wrap
		& "001"; -- Four-word burst length

begin

	-- Map ports
	nWE <= inWE;  
	iDataInput <= dataBus;
	dataBus <=
		iDataOutput when ( inWE = '0' ) else
		(others=>'Z');
	ramClk <= iThisRamClk;
	mcrDataOutput <= iThisMCRDataOutput;
	iNextRamClk <= not iThisRamClk;

	process(clk, reset) begin
		if ( reset = '1' ) then
			iThisState <= STATE_RESET;
			iThisCount <= (others=>'0');
			iThisRamClk <= '0';
			iThisMCRDataOutput <= x"DEAD";
		elsif ( clk'event and clk = '1' ) then
			iThisState <= iNextState;
			iThisCount <= iNextCount;
			iThisRamClk <= iNextRamClk;
			iThisMCRDataOutput <= iNextMCRDataOutput;
		end if;
	end process;

	-- Each state lasts 10ns @100MHz
	--
	process(iThisState, iThisCount, iDataInput, nWait, memRequest, readNotWrite,
	        iThisRamClk, mcrDataInput, mcrAddrInput, iThisMCRDataOutput) begin
		addressBus <= ADDR_HIZ;
		iDataOutput <= DATA_HIZ;
		nADV <= '1';
		nCE <= '1';
		CRE <= '0';
		inWE <= '1';
		nOE <= '1';
		iNextCount <= iThisCount;        -- by default count keeps its value
		iNextMCRDataOutput <= iThisMCRDataOutput;
		busy <= '1';
		case iThisState is

			-- 0ns: In RESET: don't come out of reset until the falling edge of ramClk, because
			-- we want there to be a rising edge halfway through the BCR write states. This
			-- ensures the BCR write works even if the RAM happens to already be in sync mode.
			when STATE_RESET =>
				iNextCount <= "0000";
				if ( iThisRamClk = '1' ) then
					-- Move on at the falling edge of iThisRamClk
					iNextState <= STATE_REQUEST_BCR_WRITE0;
				else
					-- Stay in this state whilst ramClk is high
					iNextState <= STATE_RESET;
				end if;

			-- 10ns: Assert nADV, nCE, inWE & CRE, drive BCR_INIT on addressBus
			-- RamClk is low for this state
			when STATE_REQUEST_BCR_WRITE0 =>
				nADV <= '0';                 -- tVP: nADV low for >7ns
				addressBus <= INIT_BCR;      -- tAVS: addr valid & CRE high >5ns before nADV rising
				CRE <= '1';
				nCE <= '0';                  -- tCW: low min 85ns (9 clks @100MHz)
				inWE <= '0';                 -- tWP: low min 55ns (6 clks @100MHz)
				iNextCount <= x"0";
				iNextState <= STATE_REQUEST_BCR_WRITE1;

			-- 20ns: Just in case RAM is already in sync mode, hold things stable for a ramClk rising
			-- RamClk is high for this state
			when STATE_REQUEST_BCR_WRITE1 =>
				nADV <= '0';                 -- tVP: nADV low for >7ns
				addressBus <= INIT_BCR;      -- tAVS: addr valid & CRE high >5ns before nADV rising
				CRE <= '1';
				nCE <= '0';                  -- tCW: low min 85ns (9 clks @100MHz)
				inWE <= '0';                 -- tWP: low min 55ns (6 clks @100MHz)
				iNextCount <= x"0";
				iNextState <= STATE_REQUEST_BCR_WRITE2;

			-- 30ns: Deassert nADV to clock in BCR_INIT, keep asserting nCE, inWE & CRE
			-- RamClk is low for this state
			when STATE_REQUEST_BCR_WRITE2 =>
				addressBus <= INIT_BCR;      -- tAVH: addr valid & CRE high >2ns after nADV rising
				CRE <= '1';
				nCE <= '0';                  -- tCW: low min 85ns (9 clks @100MHz)
				inWE <= '0';                 -- tWP: low min 55ns (6 clks @100MHz)
				iNextCount <= x"6";          -- Nine states = 2 + (6,5,4,3,2,1,0) = 90ns
				iNextState <= STATE_WAIT_BCR_WRITE;

			-- 30ns: 2x REQUEST states plus 7x this state gives 90ns, which meets tCW>85ns
			-- The state entered on ramClk falling edge and
			--   left on a rising edge if init iNextCount even
			--   left on a falling edge if init iNextCount odd
			when STATE_WAIT_BCR_WRITE =>
				nCE <= '0';   -- tCW: low min 85ns (9 clks @100MHz)
				inWE <= '0';  -- tWP: low min 55ns (6 clks @100MHz)
				iNextCount <= iThisCount - 1;
				if ( iThisCount = "000" ) then
					-- Last wait state before we move on
					if ( iThisRamClk = '0' ) then
						iNextState <= STATE_PREPARE_READ;      -- If the iNextCount init was odd
					else
						iNextState <= STATE_FINISH_BCR_WRITE;  -- If the iNextCount init was even
					end if;
				else
					-- Count not zero yet, so loopback...
					iNextState <= STATE_WAIT_BCR_WRITE;
				end if;

			-- OPTIONAL: ramClk was high at the end of STATE_WAIT_BCR_WRITE, so
			-- wait for ramClk rising edge before starting initial read. This state is only
			-- needed if iNextCount is initialised to an even number in STATE_REQUEST_BCR_WRITE1.
			-- Bus definitely now in synchronous mode.
			-- RamClk low during this state.
			when STATE_FINISH_BCR_WRITE =>
				iNextState <= STATE_PREPARE_READ;
			



			-- Keep nCE disabled, meeting tCBPH>8ns
			-- Bus definitely now in synchronous mode.
			-- RamClk is high during this state
			when STATE_PREPARE_READ =>
				iNextState <= STATE_REQUEST_READ;

			-- Initiate sync read of address zero
			-- RamClk has a rising edge half-way through this state
			when STATE_REQUEST_READ =>
				addressBus <= mcrAddrInput;      -- tSP: addr valid >3ns before ramClk rising
				nADV <= '0';                  -- tHD: addr valid >2ns after ramClk rising
				nCE <= '0';
				if ( iThisRamClk = '1' ) then
					iNextState <= STATE_WAIT_READ;   -- Move on
				else
					iNextState <= STATE_REQUEST_READ;  -- Hold steady after rising edge
				end if;

			-- Keep asserting nCE, assert nOE and spin whilst the RAM asserts nWait
			-- This state entered on ramClk falling edge and left on ramClk rising
			when STATE_WAIT_READ =>
				nCE <= '0';
				nOE <= '0';
				if ( nWait = '1' and iThisRamClk = '0' ) then
					-- Only proceed if nWait not asserted and ramClk is low
					-- iDataInput will be available at the end of this cycle
					iNextMCRDataOutput <= iDataInput;
					iNextState <= STATE_FINISH_READ;
				else
					-- RAM still asserts nWait, so stay in this state
					iNextState <= STATE_WAIT_READ;
				end if;

			-- RamClk high during this state
			when STATE_FINISH_READ =>
				--busy <= '0';
				nCE <= '0';
				nOE <= '0';
				iNextState <= STATE_IDLE;




			-- Deassert nCE & nOE
			when STATE_IDLE =>
				busy <= '0';
				if ( iThisRamClk = '0' and memRequest = '1' ) then
					if ( readNotWrite = '1' ) then
						iNextState <= STATE_PREPARE_READ;
					else
						iNextState <= STATE_PREPARE_WRITE;
					end if;
				else
					iNextState <= STATE_IDLE;
				end if;




			-- Keep nCE disabled, meeting tCBPH>8ns
			-- RamClk is high during this state
			when STATE_PREPARE_WRITE =>
				iNextState <= STATE_REQUEST_WRITE;

			-- Initiate sync write of address zero
			-- RamClk has a rising edge half-way through this state
			when STATE_REQUEST_WRITE =>
				addressBus <= mcrAddrInput;      -- tSP: addr valid >3ns before ramClk rising
				nADV <= '0';                  -- tHD: addr valid >2ns after ramClk rising
				nCE <= '0';
				inWE <= '0';
				if ( iThisRamClk = '1' ) then
					iNextState <= STATE_WAIT_WRITE;   -- Move on
				else
					iNextState <= STATE_REQUEST_WRITE;  -- Hold steady after rising edge
				end if;

			-- Keep asserting inWE & nCE; drive dataBus & spin whilst the RAM asserts nWait
			-- This state entered on ramClk falling edge and left on ramClk rising
			when STATE_WAIT_WRITE =>
				nCE <= '0';
				inWE <= '0';
				iDataOutput <= mcrDataInput;
				if ( nWait = '1' and iThisRamClk = '0' ) then
					-- Only proceed if nWait not asserted and ramClk is low
					-- iDataOutput will be written to RAM on the rising edge
					iNextState <= STATE_FINISH_WRITE;
				else
					-- RAM still asserts nWait, so stay in this state
					iNextState <= STATE_WAIT_WRITE;
				end if;

			-- Hold data there to meet tHD
			-- RamClk will be high for this state
			when STATE_FINISH_WRITE =>
				--busy <= '0';
				nCE <= '0';
				inWE <= '0';
				iDataOutput <= mcrDataInput;
				iNextState <= STATE_IDLE;


		end case;
	end process;
end Behavioural;
