--
-- Copyright (C) 2010 Chris McClelland
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2009 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 11.1
--  \   \         Application : xaw2vhdl
--  /   /         Filename : ClockGenerator.vhd
-- /___/   /\     Timestamp : 06/04/2010 00:04:17
-- \   \  /  \ 
--  \___\/\___\ 
--
--Command: xaw2vhdl-st C:\Users\chris\src\vhdl\test007\ipcore_dir\ClockGenerator.xaw C:\Users\chris\src\vhdl\test007\ipcore_dir\ClockGenerator
--Design Name: ClockGenerator
--Device: xc3s1200e-4fg320
--
-- Module ClockGenerator
-- Generated by Xilinx Architecture Wizard
-- Written for synthesis tool: XST

library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;
library UNISIM;
use UNISIM.Vcomponents.ALL;

entity ClockGenerator is
	port (
		CLKIN_IN        : in    std_logic;
		RST_IN          : in    std_logic;
		CLKFX_OUT       : out   std_logic;
		LOCKED_OUT      : out   std_logic;
		CLK0_OUT        : out   std_logic
	);
end ClockGenerator;

architecture BEHAVIORAL of ClockGenerator is
	signal CLKFB_IN     : std_logic;
	signal CLKIN_IBUFG  : std_logic;
	signal CLK0_BUF     : std_logic;
	signal GND_BIT      : std_logic;
begin
	GND_BIT <= '0';
	CLK0_OUT <= CLKFB_IN;
	CLKIN_IBUFG_INST : IBUFG
		port map (
			I=>CLKIN_IN,
			O=>CLKIN_IBUFG);
   
	CLK0_BUFG_INST : BUFG
		port map (
			I=>CLK0_BUF,
			O=>CLKFB_IN
		);
   
	DCM_SP_INST : DCM_SP
		generic map (
			CLK_FEEDBACK => "1X",
			CLKDV_DIVIDE => 2.0,
			CLKFX_DIVIDE => 1,
			CLKFX_MULTIPLY => 2,  -- 96MHz
			CLKIN_DIVIDE_BY_2 => FALSE,
			CLKIN_PERIOD => 20.833333333,  -- 48MHz IFCLK
			CLKOUT_PHASE_SHIFT => "NONE",
			DESKEW_ADJUST => "SYSTEM_SYNCHRONOUS",
			DFS_FREQUENCY_MODE => "LOW",
			DLL_FREQUENCY_MODE => "LOW",
			DUTY_CYCLE_CORRECTION => TRUE,
			FACTORY_JF => x"C080",
			PHASE_SHIFT => 0,
			STARTUP_WAIT => FALSE
		)
		port map (
			CLKFB=>CLKFB_IN,
			CLKIN=>CLKIN_IBUFG,
			DSSEN=>GND_BIT,
			PSCLK=>GND_BIT,
			PSEN=>GND_BIT,
			PSINCDEC=>GND_BIT,
			RST=>RST_IN,
			CLKDV=>open,
			CLKFX=>CLKFX_OUT,
			CLKFX180=>open,
			CLK0=>CLK0_BUF,
			CLK2X=>open,
			CLK2X180=>open,
			CLK90=>open,
			CLK180=>open,
			CLK270=>open,
			LOCKED=>LOCKED_OUT,
			PSDONE=>open,
			STATUS=>open
		);
   
end BEHAVIORAL;
